module Data_mem(
    input clk,
    input 
);

endmodule