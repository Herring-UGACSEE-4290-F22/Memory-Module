module RAM(
    /*
    * ???
    */
);

endmodule